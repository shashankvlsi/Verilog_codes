module datatypes();
reg a;
wire b;
wor c;
wand d;
integer e;
real f;
tri g;
tri0 h;
tri1 i;
supply0 j;
supply1 k;
time l;
initial
#1 $display("a=%b b=%b c=%b d=%b e=%b f=%b g=%b h=%b i=%b j=%b k=%b l=%b",a,b,c,d,e,f,g,h,i,j,k,l);
endmodule
