module operator();
reg[3:0] a,b;
reg[16:0]y;
reg s;
initial
        begin

a=11;b=6;#10;
y=a+b;
$display("Airthmatic Operators");
$display("add y=%0d",y);
y=a-b;
$display("sub y=%0d",y);
y=a*b;
$display("multi y=%0d",y);
y=a/b;
$display("divide y=%0d",y);
y=a%b;
$display("mod y=%0d",y);
$display("--------------------------------------------------------------------------------------------------------");
$display("Logical Operators");
y=a&&b;
$display("and a=%b b=%b y=%0b",a,b,y);
y=a||b;
$display("or a=%b b=%b y=%0b",a,b,y);
y=!a;
$display("not a=%b b=%b y=%0b",a,b,y);
$display("--------------------------------------------------------------------------------------------------------");
$display("Bitwise Operators");
y=a&b;
$display("and a=%b b=%b y=%0b",a,b,y);
y=a|b;
$display("or a=%b b=%b y=%0b",a,b,y);
y=~a;
$display("not a=%b b=%b y=%0b",a,b,y);
y=~(a&b);
$display("nand a=%b b=%b y=%0b",a,b,y);
y=~(a|b);
$display("nor a=%b b=%b y=%0b",a,b,y);
y=a^b;
$display("xor a=%b b=%b y=%0b",a,b,y);
y=a~^b;
$display("xnor a=%b b=%b y=%0b",a,b,y);
$display("--------------------------------------------------------------------------------------------------------");
$display("Relational Operator");
y=a<b;
$display("less a=%b b=%b y=%0b",a,b,y);
y=a>b;
$display("greater a=%b b=%b y=%0b",a,b,y);
y=a<=b;
$display("LE a=%b b=%b y=%0b",a,b,y);
y=a>=b;
$display("GE a=%b b=%b y=%0b",a,b,y);
$display("--------------------------------------------------------------------------------------------------------");
$display("Equality Operator");
y=a==b;
$display("E a=%b b=%b y=%0b",a,b,y);
y=a!=b;
$display("NE a=%b b=%b y=%0b",a,b,y);
y=a===b;
$display("CE a=%b b=%b y=%0b",a,b,y);
y=a!==b;
$display("CNE a=%b b=%b y=%0b",a,b,y);
$display("--------------------------------------------------------------------------------------------------------");
$display("Reductional Operators");
y=&b;
$display("and a=%b b=%b y=%0b",a,b,y);
y=|b;
$display("or a=%b b=%b y=%0b",a,b,y);
y=~a;
$display("not a=%b b=%b y=%0b",a,b,y);
y=~(&b);
$display("nand a=%b b=%b y=%0b",a,b,y);
y=~(|b);
$display("nor a=%b b=%b y=%0b",a,b,y);
y=a^b;
$display("xor a=%b b=%b y=%0b",a,b,y);
y=~^b;
$display("xnor a=%b b=%b y=%0b",a,b,y);
$display("--------------------------------------------------------------------------------------------------------");
$display("Shifting Operator");
y=b<<2;
$display("lls a=%b b=%b y=%0b",a,b,y);
y=b>>2;
$display("lrs a=%b b=%b y=%0b",a,b,y);
y=a<<<2;
$display("als a=%b b=%b y=%0b",a,b,y);
y=a>>>2;
$display("ars a=%b b=%b y=%0b",a,b,y);
$display("--------------------------------------------------------------------------------------------------------");
$display("Conditional Operator");
s=1;
y=s?a:b;
$display("CO a=%b b=%b s=%b y=%0b",a,b,s,y);
s=0;
y=s?a:b;
$display("CO a=%b b=%b s=%b y=%0b",a,b,s,y);
$display("--------------------------------------------------------------------------------------------------------");
$display("Concatenation AND Replication");
y={a,b,a,b};
$display("concatenation a=%b b=%b y=%0b",a,b,y);
y={4{a}};
$display("Replication a=%b b=%b y=%0b",a,b,y);

        end

endmodule
